push int8(100) ; d
push int8(108) ; l
push int8(114) ; r
push int8(111) ; o
push int8(87) ; W
push int8(32) ; SPACE
push int8(111) ; o
push int8(108) ; l
push int8(108) ; l
push int8(101) ; e
push int8(72) ; H
print
pop
print
pop
print
pop
print
pop
print
pop
print
pop
print
pop
print
pop
print
pop
print
pop
print
pop
exit