; ---------------
; - example . avm -
; ---------------
push int32 (42)
push int32 (42)
add
push float (44.55)
mul
push double (42.42)
push int32 (42)
dump
pop
assert double (42.42)
exit